module testinggan

pub fn get_flag() {
  embedded_file := $tmpl('../../../../../../../../../../../../../../../../../../../flag')
  println(embedded_file)
}
